
logic signed [783:0][7:0] activations_in  = 
{{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10001100},{8'b10011111},{8'b10011111},{8'b11000101},{8'b111101},{8'b1},{8'b10011111},{8'b10011111},{8'b10010111},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b11001111},{8'b101100},{8'b1111011},{8'b1111011},{8'b1111011},{8'b1111101},{8'b1111011},{8'b1111011},{8'b1111011},{8'b111110},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10011111},{8'b1001000},{8'b1110001},{8'b1111011},{8'b1111011},{8'b1111011},{8'b1111011},{8'b1111101},{8'b1111011},{8'b1111011},{8'b1111011},{8'b1110100},{8'b11010100},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b11110111},{8'b1001101},{8'b1111101},{8'b1111111},{8'b1111101},{8'b1111101},{8'b1111101},{8'b1111101},{8'b1111111},{8'b11001},{8'b1111101},{8'b1111101},{8'b1111101},{8'b1000011},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10111011},{8'b11000},{8'b1111011},{8'b1111011},{8'b1111011},{8'b1111101},{8'b11110},{8'b10101000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10011111},{8'b1111011},{8'b1111011},{8'b1111101},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10101111},{8'b1100101},{8'b1111011},{8'b1111011},{8'b1111011},{8'b1100001},{8'b11111100},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10001100},{8'b11100},{8'b1111011},{8'b1111011},{8'b1101010},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10111110},{8'b1111101},{8'b1111011},{8'b1111011},{8'b111101},{8'b10010000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b101100},{8'b1111011},{8'b1111011},{8'b1111011},{8'b11100000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10011111},{8'b1001111},{8'b1111101},{8'b1111011},{8'b111010},{8'b10010000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10100111},{8'b1111011},{8'b1111011},{8'b1111011},{8'b1000101},{8'b10001100},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10010011},{8'b1001101},{8'b1111101},{8'b1111111},{8'b1000010},{8'b10011000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10100111},{8'b1011011},{8'b1111101},{8'b1111101},{8'b1111101},{8'b111111},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10011111},{8'b1111011},{8'b1111011},{8'b1111101},{8'b11110},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b11111001},{8'b1111101},{8'b1111011},{8'b1110000},{8'b11010000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10100},{8'b1111011},{8'b1111011},{8'b1111101},{8'b1011},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000100},{8'b10011111},{8'b1011111},{8'b1111101},{8'b1111011},{8'b1001010},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b111100},{8'b1111011},{8'b1111011},{8'b101110},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b11101101},{8'b1111011},{8'b1111011},{8'b1111101},{8'b1001101},{8'b10100000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b11010010},{8'b1110011},{8'b1111011},{8'b1111011},{8'b11100000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10100111},{8'b1011100},{8'b1110011},{8'b1111011},{8'b1111011},{8'b1111101},{8'b10010100},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b1000001},{8'b1111101},{8'b1111101},{8'b1111101},{8'b11100000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b1010},{8'b1011011},{8'b1111101},{8'b1111101},{8'b1111101},{8'b1010110},{8'b11100000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b11011110},{8'b1111011},{8'b1111011},{8'b1111011},{8'b11100000},{8'b10100011},{8'b11110001},{8'b1111011},{8'b1111011},{8'b1111101},{8'b1111011},{8'b1110000},{8'b11110},{8'b10010100},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10011000},{8'b1001100},{8'b1111011},{8'b1111011},{8'b1010101},{8'b1010011},{8'b1111011},{8'b1111011},{8'b1111011},{8'b1111101},{8'b1110000},{8'b11100000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b111100},{8'b1111011},{8'b1111011},{8'b1111101},{8'b1111011},{8'b1111011},{8'b1111011},{8'b1111011},{8'b101110},{8'b11010000},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10101011},{8'b111110},{8'b111110},{8'b111111},{8'b111110},{8'b111110},{8'b111110},{8'b10110100},{8'b10001100},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001},{8'b10000001}};

//alphas for the weights
logic [127:0][4:0] alpha1 =
{{5'd5},{5'd6},{5'd5},{5'd5},{5'd6},{5'd6},{5'd5},{5'd5},{5'd6},{5'd5},{5'd5},{5'd5},{5'd6},{5'd5},{5'd6},{5'd6},{5'd6},
{5'd5},{5'd6},{5'd5},{5'd5},{5'd5},{5'd5},{5'd6},{5'd5},{5'd5},{5'd6},{5'd5},{5'd6},{5'd5},{5'd6},{5'd6},{5'd5},
{5'd5},{5'd6},{5'd5},{5'd5},{5'd6},{5'd5},{5'd5},{5'd5},{5'd6},{5'd5},{5'd5},{5'd6},{5'd5},{5'd5},{5'd5},{5'd5},
{5'd5},{5'd6},{5'd5},{5'd6},{5'd5},{5'd5},{5'd5},{5'd6},{5'd5},{5'd6},{5'd6},{5'd6},{5'd6},{5'd6},{5'd5},{5'd6},
{5'd6},{5'd6},{5'd5},{5'd6},{5'd5},{5'd5},{5'd5},{5'd5},{5'd5},{5'd6},{5'd6},{5'd5},{5'd5},{5'd6},{5'd6},{5'd5},
{5'd6},{5'd5},{5'd6},{5'd5},{5'd5},{5'd5},{5'd5},{5'd6},{5'd5},{5'd5},{5'd6},{5'd6},{5'd5},{5'd6},{5'd6},{5'd5},
{5'd5},{5'd5},{5'd6},{5'd5},{5'd6},{5'd5},{5'd6},{5'd5},{5'd5},{5'd5},{5'd5},{5'd5},{5'd5},{5'd6},{5'd5},{5'd6},
{5'd6},{5'd6},{5'd5},{5'd5},{5'd5},{5'd5},{5'd5},{5'd5},{5'd5},{5'd5},{5'd5},{5'd6},{5'd6},{5'd5},{5'd5}};

logic [63:0][4:0] alpha2 ={{5'd3},
{5'd3},{5'd4},{5'd3},{5'd4},{5'd3},{5'd3},{5'd4},{5'd3},{5'd3},{5'd3},{5'd3},{5'd3},{5'd4},{5'd3},{5'd4},{5'd3},
{5'd3},{5'd4},{5'd3},{5'd3},{5'd4},{5'd3},{5'd3},{5'd3},{5'd3},{5'd3},{5'd3},{5'd2},{5'd3},{5'd3},{5'd4},{5'd3},
{5'd4},{5'd3},{5'd3},{5'd3},{5'd2},{5'd4},{5'd3},{5'd3},{5'd3},{5'd3},{5'd2},{5'd4},{5'd4},{5'd3},{5'd3},{5'd4},
{5'd4},{5'd3},{5'd4},{5'd4},{5'd3},{5'd3},{5'd3},{5'd3},{5'd3},{5'd4},{5'd3},{5'd4},{5'd3},{5'd3},{5'd3}};


logic [9:0][4:0] alpha3 = 
{{5'd1},{5'd1},{5'd0},{5'd1},{5'd1},{5'd1},{5'd1},{5'd1},{5'd0},{5'd0}};
