logic  [127:0] [783:0] input_weights= 
{{784'b0111001011011101011110111001001110011011001010011111011110110110110011010011000100101100100100110100100011000111111101000110000011010000100011101000111010000000111001010010111111101100010000111011111011111111100000011101001010100011111111000111111111101111101111111001111010110111101011010010110011001010111001001100001000001100000001111001000000000000011000000011110010100000000001001001101111100000001000001100001111100011100001100000011100110011000000000010000111001101111001111011010000011010001111101111000100001110011000000011001010001011111100000101110011100010110111100001000011101010100000011111010000111111011100001101111101101011011111000101101010110001111111011110111000001111101111101101110111001001101111101011011111101100101000001000110111001011111111001000000011111101},
{784'b0100101011001101100100001011101100101011101111011100001101100101010000011001110101010110101100001010111001111111010011010000011110010111001100110000000001010000101100111110111000010110000001010010111111001100101010111001010100110000111000011111010001001110111000000011001111100011110010011000001111110111000000001101111110111011111011111011111111111111001111100111110001111111100101000111001011101110000000001100000101000001101111100001110010000011010110011100100000010101101010000100010001010001001010111000000101101110000100000010011000000000110000111001000110011000000001100000000011110101000011101111001001000101111001000100101010010100010111110111010101000001011111110100101101110110010011100111101001001110001100011010110100110010011111001111111111111011111010011010110111011110},
{784'b0110011101001110110111111101110111110111011111110011011111101011111110010011101011110110111101000000011111111011011101110000000010001101110010001100000000010101000111011100110000011010010010111110101001000000001111001111110010100000000011111101111011001001100000000111010111101111111010000000111011110111111111110000000111110111000101110000000000111111001000000011111010000111111000001000011001000000001111011001110000001110000000001011111010000101111101000001110111100000000110111000000001111110000000010011000000010111111000000111111111101000111111100000000111100010011000111000000000100010001000001001000000001101111110100111111100000000000011100111111111100000000010111111111111111100000000010111001010111111100000111101011011010111111111111111011101010000101100110101100111101001},
{784'b1001001000110011110011001111101011110001001100110101111111101011001111010010101001101111110001111101001111101011110011001000000000010110110111011010000100000000000011100001101011100000001001101000011011111111111011001100000110101111111100000111000000101011111111111001110100000010111101111000001111000000001110111010000000111111100000100111100000000111111010000111101000000001011111110101111110011000011111111111010010111001000011111111111111110010110100011111111110110010001010011000000111111010010100111011000000000110001101000000011110000000000000000000011111111000000000000000010011010101111000100000000000000010101101111110010000000001101011101111101111000000000011101000111101100000000000101100110011111101110011011110111110110011111011111001010111101111111000111110011111101011},
{784'b1110110111011010000101101011111000000101000100010101011111001111101110111001010010111110011010111101101001100111010011110000110110001101111101000111011101010110000101101010011000000111010011100011111011011010110110101100101110111011001101111000001101100011101000111110110000110110110010011010111001001111000011010111000011100000011110010011011101011100110110111111001001100011100010001111111010110100000111010101010011101111000001111001001110011000001111101111100011111100111010010111011100001111000111110110011011111101110001010011110111000111100001000100011110011000111110010000011000011000111101011001000000100101001110110111110000000010001011101011010001100000010111110011001101111110000101011101101100101101011100001010110101011111000000000101001100000110111111001010010010101000},
{784'b1000010001101110101000101101001100000001111010101001000001100100110110101100100110010011001101011000101101011100111011011110111011111101001001111010110001001001111101100001111011101010101010000101010111011100000101100010100110110110101100011111011010111010111000000000001010101101010011000000000010111001000000101000000000001010010000100111000100110010111010000000111001000001000111110001010101000000101100011111111101011110001111010111011101100011110010111001111100110111100110010001100110110110111111000001110001111110111101000111111000010011111110010110010010100001000001100110100010100010000000101111001110000111010011111010110100001101101000101010001100110100101000010000011100100010111000000101111100011111111101110111100100101100100001101111000001011000110100010011101110110011},
{784'b1111000010010111111011000011110111000101101100101110100101110111010010110001110100101011111110111111111000011001111111000101111101101011100011101111010111111010101111010101001001111111000000001011110110000111111000000000000111000000111110000000000001011001101111111101000000001110111000111111111111000101111001100011101001111111000011111000001111011011011011000100100010111011101010001000010011000011001110000000011010111101100100110100000000011011010000000001100001111010000111011000000000100101000011011001000100000001111000000010000000011000001111001111110110000100010101011101001110111101001111111000000101111011010111110111010000111011001110111010101100100110111011111100100010100000010010111111111011110011000111100111000111000110010111101101110111010101101100010011001101001001},
{784'b0110001010000010110000101111001101100111010110010001010011110101101101110001101101001011000011111000010000010000100010100110101011001010111010011111100011000010011100011110101101100011100011011001101100001001001010001001011110111001011001110011011100111000001000100010111111110110001001011100011011111111110011101011000001100111111110011010011000001110100001111010111100010000111001000000111001111011000011110000001101010100101100000111100000001100101111110000001110000010111100101111000100011100000001101111111111010011100000011100000101111101001110000011000011010011111111111000000010010101111010111111000000111000001011111111110000000011101010010001111111000000010001000010100111101000000100100111010000000101000001000011111000010011000111100111011101100000110000001110101000100000},
{784'b1110110001011010010101111100100101010010111010100011110111110111111110101000101101110001111011111111110000110101001001011110111111000001110001110111101001011000000001111111010010011110101000000010011000000010101100010000001001100000001110100111011000110101110000110111111010000101000010100000111111101000011101000000000001011011110000000111100001000011111111100010110000000000011111010001100101110000100010100010110001110000101111011101100000101111101010100110011011110000111110011010010000100000101011110011010110010001110111101100011100000110111101101111110001100110111010101011111110101011101110100100011110111110110110000010000010001000011100110110000000000011010111000001001101000000010100011010110101011000110000101010000101101101101111100101111001111111000110101000100100000101},
{784'b1101000111011001001011000011100110101101111100110001000001110100001111000010010011101000010101100101111010100001100110110010010110110100001111011011011000000001101001110110111100100000001101000010111001010010000011111100000100101000011110001111111000111001010111111001111111110110001001011111000111101110000100111110111000011110000000101001101111000001101011100111101101111000000001001111111100110111000000000000000110111001100000000001000010010101111011100000000000001101101110111001100100000000010111100101111101111000001111101111110111111111110011111111000110111011111111000110101110000001010111111000001011100111101011101100001001111111000101101111000010000100101000100110111000000000011011111010100001001100111101000110000111000100000011010000001101011101011001100110001010111101},
{784'b1001100110101100101110010010100111101111111010011000001011000100101000000000000000111100010101000101000010010010110111001000110100000100100001001101101111111011010110000001000111011110101101110011011110001110010000001110011001100100111000110001111101111001000101111111110010010000111000110111111111110101010010110010000000111100000000001000001101001111100000000110100000110000111101100011001000011101110111001110011000111110100111111000010110010110001010111110000010111111010010011111111000000000111110000000111111000000100011110000010011111000000000011111110010001111100001100010111101100101101110001001100111110110001001111011101001111111010111010001110100100011111001001001000010000000000011001001010110010000000000001001011010010110111100110010000001110000101100111111010101100100},
{784'b1101111111110111011100110100100010101011111111010001100000110110110110010011111101011111111000100000000001110100101011100001001110101000101000111100100011111110001111111011111011001010110000101000111111111100100000000010101001000100110001111001011100110100011101110011110010111010111101110111101110011111010110111010111010100011111110110110100111101010011111110110110001111111111100111111001110011001111111111100011100010011100001111111100000001011001100000001111110000000110101100000000001000000011000111010010000000000000000100111000110000000000000000101000110000110000001000010000001001110111110111101000010110000110001111111011000000111111110111001101111100101000000011101100111100000000011011110001000100100110000011101100100011111101010100100010010111110101101001100110000101001},
{784'b1101101110100011101011000101111001001110000101000101100101000010010111101111110101000000011100110111000011111101111000011100010111000101111111011111001000010000011000111001000100010011000000110010111000000001001110000111111111011000100100100000010111110101001010000111000011001001111110010101010100000101011100000000101000011011000100100100100011000100000000000000110100000010111011100001000111100100111011111000000010101111000111111100110000001011011000100111001001000000010111011010011101111110000111101000011111101111110111011110001111010011111111101011001001110001111111111111000111110110110011111110111111110101111101011011101110111000011011100100000010010001001111011100000100011010011101001001010011100100011001011100000011110000111111111100000001010100011111101110111000001011},
{784'b1110100010101000110110010001100010100000011100000101010001010011011100110010101010011101010010110001111011000000010010001110111110011110100011011111011111111001111110111110011111111111000011110110110001111111111000000001101110110111111110000000000111101101101111010000011001110110010110010100000011101111111010000000001000011111001101001000001111101001110110100110001011101110000111001100000000000101100000010011000110100010010100000010000101000010110110001100111100000010001100101001010111100000001100010000101100011100000001010011011000110100000011101110010010001001101000011111110100010110011111010011111111100111101001111111011111111101001101011000110111111111100100010000000001111111111110101100110000110000000101000000010110110000000000000001110100100000010000110100110000011100},
{784'b0001110001001000010101011101000101011010001101010001010110001011101010110011100010000001001000011110100000010110111110101111100111100000111000000101111111111000100001100000110010101111111110000001111100000101110111111010000100000010101001110110110110111001001001101111100100100010100101111111011110010110001010111111111100110101101100100001111111000010100110000111000110000000011101101110111000111010100011011010000000001001001000001011110001101011100010001010010100000100100001101101000011000100011100010110111101010000001010110110100100000011100001011011000100010100110011100011011101110001110011001001000001111111000100011000001010011110111011111011011110011010101111000001110100010001010110111110001111001010000110011110111100001111111101111110111000111111100101100001100111111010},
{784'b0011011111001110111111010110001101100000000100110110000100111010100011100111111011011111110100000101111001001111110100110111100011100000010101111101111111110010100110100001101101101111001100101011001001001110111110000101011011110001100101111001110010111011101100000111101111001001111110010100001111001010010011111001011111110111011011011110111010111100100100101110101101111110100000001011100010111111010000000001111001111100010110000000000010011111110011110000000000011011101111100011101010000110010101111110110000100000011110010001011000010000100000101010000010010000000100000100011000100011000000000001000010001010000110101011010101000001011001110110010011110001000011110001111100100111100010010110111010111111110011010011100101001001100010100010110101100010111000010000110110111111},
{784'b1010111111011111000011101101111101110101111110011101111010111111101001100111101100111001101001100100001100101011100110000000000000001011011011111001000011100100111001111100110010111111110110011111011100000100111111010100100100100000000001011000011011100100001000011111001000011110101100001011011000000010111111111010001101111100000011111010111010001111111000000111110111000000010111111000010001100000010001000000000001101100010110110000110000000111011110111011000011111000111111101111100011001111100000111011101111111011101110000000111111101101101010010100100100110000110100010110000011000100001000001001101101101011101111000111000010001001000010100110000100000000111111111011101000000000111011110101000111010111100101111110101101100011101100110111000011100111011111001101101111111100},
{784'b0000001111010000001101000110000110101111100111011000001001000000000010100010000111101000100000010001010000001101100011111011110101110000100010110001111111011000101111011010111111111111110001001110010111111111111111100110110100011111111101111011001111010010111111111111011001001111010010111111111101101000011111110110111110111110000011100001111111111111101100000111011110000101111111110000010010010000000001111110000001110111000000000111110001010010111110000000000111000001010110110000000000111100000111110001101000000011110110110010110110101000010111000101100100010011000001001010000000101100101110101110101001000110100111011111001001110000101100110111001011101111110110110100101111111011010111100100101111111111111000111100101000001000110100101011111000001000010101001100110000111000},
{784'b0110000101010010010101101010000010101000101100011100100100011001000110111111101001100000110110111111011111101101100110100111110101001010000000101011111011011100001000010000011001000001000000100000010001110111011100100000100010111101011111111001010000101000111111111011011001000000001100111010001010011111001100101001000000111111111110010011100001000010111011111100111110100010001001101101101001000000100000010111010111110100011100000101010111111000000111100000010000000010101010000001000010000001111110010100010010001111001000111000000001010010111100111111010000011101101110000001101011110010011101001010000010001001000100111111000100000000110001001011100011001100000100000001010100100100100001100011001010111111111101111101100010111101111111111111000111001010101001101001000011001010},
{784'b1000100010011011110110010011010110001011010001010000100001011000000000010010000010101110111000100000000000110011111101011101010010011011100110010111010111111111111100010100001110111111111110110001011011111111111111111111100100010011111111111110101000000001101111110000000000000001000010100100000000010010000101100100100000000000000000100100000000000000001111000000101110000101101111100011111011010011110111111100000001101101110101110111110000010011000110111111111111000010111010100000001111111100101111000110110000000011101011100110001100100000000011001101101011001001000000000001111011011111100100010000000111110010000111111111111101111111111000001011010111111111110111010000110011111000101100101010111101000110000000000010010011010100010000000111011101111101011100001101000001111000},
{784'b1100011010011111111111110111100001100011011110011101100110111011001001010000010001010111010001000001111110000111011110010000001000111001011101110001000100001111010110001000100000000011100111111111101100001000111100111100000000000001111110011110111111010101001111110000000111110011110010111110000001111110111111111111000000011110001000111101100000000001101101001111011000000000110011111001111011100000000111111000010000000000100001111111000001001111101111111111111100000101101110110001111111110111000101010111111100000011111100001011001011110000000011000010110110011111001000010010101101100010111000001101111000011010111000111001001100101101011110001110000001011101101101101101011100101010110100001010011111111110010011001000101101101100000100001100000010111010111100000110111011101001},
{784'b1110000110110000000100011001110010101110110101011111001110111100010000110000100000010011100000000000101000001011000101000010110000100000011110010011111000110010111011000101100111100101111100010100101101111010011111111000100001001100101100111111010001110110001010000111111100110101001000100100000111110111110101111100000000011110000011000100111101100000100010000101100111111110000010000010001100110101110000011111011100011111111100000000110011000010110101110000000111111010111010110110000000111110111111001111111100000011011100000001000111000000011111110100000101000110100001111101000000001010101100001011111110000101011111010100000001111011010111011111110000000100010011011011111101100000000001000010101101011100101000000110110000111111111101011101011011011110111010110000000100000010},
{784'b0000111000100001110110010000010011100111000011110000010000101010110000100001000111000111100000000011000110010100000110000100101111111001010100100000001001011111111100000010000100000101111111111100100100111111110011111111010001010010100110100111111111110001001001110000111111111110100111111110000011110011110110011111110000011111100001010001001100000111100011100010000011010000001101000000000100111100011111100100010010011100110010111101001100001000010000100011110001100100010111000110111110010010000011100000011101111100000010001111111011111111001100110000011001001110101100000101111101111000011111011011100101111010010111111100111011100011100010101011111110111010000110111011110001000000010100100000010100101000110111111110011100010010011011111111110110110010000110100001000011000000},
{784'b1111101010000001111110110011001011101110010111111001010000011100100010100100100000101010100100000000000100001010010110110000000011010110101100101101000001110111011001101110001110011000010111010111110111100010101101110111010000111111111010011011001110010110111110000000111111100111100110010010111100110111000101000101011111010101001011010011001011111110111111010110001110101111100111101100110110111101110100111101100001101111010101111000111010000100011100001100101101000001000111001001011011101001000000101010010000001101000001000000111001110000000000000000000101111011000000000110011001011100000000000000010101000101110000110010111111011100100110110110011111111111010011000111011100110110010001000011110001101111001110110000101011110100000101000110001110111110111110001110111111111101},
{784'b1001000010000000011101011010100001000101111001110011110010011100100111110101101111010111000110001001110101110000001000001000010001111000111010100000110110000110010010101010001000100000000010000001100100001000000000000000100001100111010000000000111100111111001111110000011111101110010111111111100011110111011111111111111111111111111111010111111111111111111111111001110101011111111111011111000100111111011111111111111000000011110011111111111101101101110010111111111111101011001101100111111111111110000001011110011111111111101000001100111111011111111000000000000101000000101000000001000010010000001100000000000000000110010000000000000000001101000111110000100010000001010111100011010000000000000110110011010011100000001001001000101000000001010000000011100100101101100111011000100111100010},
{784'b0011000001001100000010101101010100101101001010010111000111001110100000101101111000010000010111000101110000000110011000000010101111111100100010110010001000111111111100100111001100000001111111111010100000101001100111111111100000000010110100000111111111001000001011110000011111111101100000111100000001111111100010000010010000001111101101111000000000100001110110000011001110110100000111110000001010000111010001111100000010100010101100011101100000000011000001100010101101010000011010000101111100001000000111000010011111110011000000011000011101111111001010101011100010111111111100001011111101011100001111111110010101110011001010111111110001001111001100110011111111100001100111001110001011111111101100100110010000000011010000001000100010100110110011001001001100100001010111111001001010010101},
{784'b1110011111110011011110000000110111101010100010101111001010110011110111111110000111101111000011000010001111100001011011110010001001000011111011101101001000000011001001111101000011000000101100010110010000001000000000000000011010010000000000000000000001011001001000001100000010100010100000111111100000010101111110000111111111111111000101110001111111111111001111110100011011111111111111111111001011111111010001111001101011111101001011000011110100100111011110101101101000000000001010011111000110111011110010100110011001101101011010000111110110110101000111100101100000000000000000101101010000010100000000000000001111101111011010000000000000011111011010011000000010001111111111101111010001000000011111111111110110000111111000110101110110100101110111111111011110011110101110001010010001111101},
{784'b0001101011001000101111011101111111001100000101010110110011110110100101000000000000101111111000010000000000000111100110001000000000000000111111110100000000000000000001001111001000100000000000100100111100000000000000001111101010110000000100011111111101001011100000011111111111101111011100010111111111111111111010000011011111111011011001110100101111111011000000000101001100111111001000000000010011111111111110001110000110111101101111111001111001000011010011111101111111110001111101111111101111111101000101111100111111110100101111001101111011110000000110000101110000110110000000001010100101101101000000000000000000011011011110000000000000000011111111011100001000000001001111111010111110110000011111110111111000001000000001010101010100001010101011111010111001110011110111111011111101111011},
{784'b1001111111100000110101010010010000100101100100110001111111000101011011001001011110001110010101010111001110111000101110001110110011101111100101000101000000010011111100011100101100111001100010111010101010110101111111011000111110010111101110110001000000101010010100001000000000000011101111001010001110001100000010000101110011111100011100000001001011110111110111111000110001110100001110011111010000001011110000111011011111100111111111100111010111000011110010011111001110010001011100000011111111110000000001010101101001001110100010001000100010100001101101011101001011001000001011000101000010011001100010001001111111101011110111010111000100001100010010110100000000001011000011001111010100001000100100001011100001001101001111000110010100000000011111111101001101011110000011011011000001000100},
{784'b1100000101110000101001000011110001000000001010011010100011000011000100100001011000000100111001101011100101000000100101001111111000110010000010011001111011000010000100000111011111110100000010111110111010111111101001000110101000101111110001111110101100100011111111000011111110000011010111111100001111111110000010010111100000011000100100010010111111000000000001110101101110111110000000000001110100101111111100000011111010011001001111110010000111110100000000010111011000101111010001110100001111100011110101100011000000101100001111010010001110001101111100111110100000011111110110101000111111000101000101001011001111110000000110000000001111111010001000001111111101001111110101101000110101110011000101000000000100001101111000010001101010001101100111000010000001100011010100010100000101100100},
{784'b0011000000011000111100101100110100100000001100010101011001111110100011111000010111101110110011110010000101011000000000110110011010011000010101101111100000110000000000011101011000010111011101000001000111010111101111111010000010011110111011111111111100010111111011110111111111100011011111111011111111111110000110010100000001110111111000010110101000000011101101111101010000000000001100000010110001001001100010011111110111001100000010100111111110111001010011000001001010110110100110000101110001101000111111101101010000000010110101011010110100010000000001111001110110110011110001010011010001100101011110101010000000001001011110111010001100000001111001010010010001001011001101101001111111011100010111011001111100101111000000001111001110110010000110010100111011001010101000000111101001101101},
{784'b1100001101010011011111110100110011001110010010111101011011111111010000001011100100111111101011000000000101011111011110000000010000111111111110110000001100001100100111111110010001001000001110111000110011010100000110111111110111010011101000000011111111001100001100110001000001011001111111101111011110000000111011010100111111111011000011111010010011011101111010000010000000000101100110001000011111110010001100010111000001000010100000100111000101000111110011011100011010101000010110110100100111111000010010011010010111001110000011101111011101100000010111100000111100100001000000000100001001010100000000010010011101000101011010110101100011111100111110111010011001111101110101100111110001010010110100010011011011000100101010000011100101000000010000000000110100010111011011100101000010111111},
{784'b0101010101111000011001111011100010100011110010001011101111011001110100111110001000001000111001101000000000000011001110010000000000000100011111101000000101000000000010100011010000011111111000001000111110001110111110101100001111111111011111111101101110110010011111111111110100000110111101111111111111011001011111011111000001111110001111101100101000000001101100000011001100000000000011010100011000100000000000111110010001100000000000000011000001000110000001001100111100000101101100010011111111110000000011110101101110111110000110101111111101010101111010100011101001110000111100101000101111111111111011101000000110001111110011101100001000101011110101000010000010000000110101101101011010000000001111111101100011110000101101111110101011100101011110111111010111111111001111111100110110001001},
{784'b1111001110011101011110011101110101010010110011010101100011000101010001001001111110100101001110001000001001101101011011001100111111011111011110001101101011111111011010111001111110001000000000111011011111111000000000000001111110000110000100000001010101110000100000000000000011001100010100000000000001110000110010001000000011100101001011001110000011111110000001101100011100111111111000000111110101010000111111110100001111000001101111111110000110011000111101101101011100111011110000010111100110001101110110100011011011111100101001110110010101111111111111001110001010010111111111101111111100001111011111111111010001100011111101000011111110011110101111101000001011111001010011100110000000000000000100000111011100000000000000000000001010000010000000000000101101110110100000101010110000000100},
{784'b1100111110100101111110010000100111101011111010110010010010001110111010010010110011000111001010100101110010100111100000000000000110110101001110011010000100101111111011010110010000011101100101010000111001000001011100111111101011100110010011010110000100001101001101111011111010101001011010100111100000010101000101011111111111100000101110101000011111111110011111111100100111111111111100100011010110110111111101100000000000101110010111111000000000111100100011110111000000000101101111101110111100000000001110000100010111100000000111110111011001011110000000011111100100010000101110000111110101110010001001000000111111101100010000011011111111100110001011000000110111011111110001111011000101001111101011100001100100101000100001001001101000101110001011011001011010001010010011001001100100000011},
{784'b0101000100101010000101001100101100100011110110001000010000000001001101100000010100001111001001110100110101110010100001100100000011101000100101111010100100100001111110111000100011001100000011111001111000011110010000110011100100111110110100011111110110111100000100000111111111010000111101110111110000001111001110011110010000000000001000001001111001000000000010111101010100100100000000101011111000001111111111111110000101000001111111111111101000011010101000111111111110000010011100000000111111110110101000101000000001111000111110011010000000000000000101111110101000100100000000010111110100111010000000000110101111110101101010111001000011000110101001010011111101110011101101011000010101111111001000110010000010101001110001100111100101011010101101011000001000010101011111101001101101001001},
{784'b0000011100111010001010110100111101011000100110110001000101111011111010100000001010010010110111111011110110001100000011111111111001011000001100111110111110001000000001000011110101000000101000000101011011011101110111010000001101111111111000111110000000111101111100001111111110000000000111100000000111111110000000101100101100001111110001110110101001100000111111111110110110001111000111111111101011111111010000111111110100011101111010100011111111110111000011110000100111111111010011010111100011011111111010001001000110011111111110000000011011000100011111001000110110001000000001000000100101110010010010000000000000000011000100011011000000000000001001110000000100000000001011100111111100110100011010110001000011010010101111111110000000000101100000001011100001010011100110011010010001001001},
{784'b0111010110100101000110100110100101010111110000010010000111001111110110101111000000110010011111001011001100100111011100101001011101001010000010111011111001101111011010110000010110001000010100100100010100001111001001110011011111001111111011101101111100111101101001100110111110111110101000111111111111011110100110000000110111101101101010000010001101001111110001011001110100000110101001011001011110000100001101110111001000100101110101011101101011110011100010111000111111100111010100111011001111011100100011111101110010110111010000111100100000001010011000000110011001111111001100000000101000110111011101001001000110001001100111111110110111000100011001101000000010111000000011001010000000010001110000111101011101100001001010100011001010011101010100011101000110111100110010011101101111000100},
{784'b0100100110111101011010011000111000111100100111001101010111111001001010001011011111000011111100010000000100000111000101011111010000010011111111100011001110000000010010110101111010000000001101000011110010100000000000100000000110000000100000000010010001011100011101111000111110000010000111111111110111000100101111101111111110001111011000011011111111111001111101110001100111111111000011111111010100011111111000001111111111111111111111100001111111110001010101110000000110111111110011000111000000010000011010011110000000000000000000100100100000000000010010000001000001110100000010001010001000111110000000010001000000000100011100001100000000100000001101110000100000001101110010111000110010000000101111110111000011000010110001011011100000110011010011110001101010011111100100110100010101001000},
{784'b1110001111110001000000101101001010011110000001100101001000000011001011010110010010001100000010111001110111111101000111101110010101011011010101000111101100011111011110010000000000000000100111010011000100101000000011111010010010010101101000001101010001000010111110000001100110000001101010011111100011110000000000001011111110000111001011000011111111111000101100000001100011111111110000000010001100001111111000110000000000001100111110000000000011011011111001110000011010000010010101010100000001111111010111001010010000001111111111100001111011100000111011111101110000110100000111101111111000011011010000101110111111111000011010000000011111111111011010100001000000111101101100000010111100000011010101010001111011111100000001000110101011100100000110111111100100100111101101101110010000100000},
{784'b1011000010101011100110000111001000100110110001100100001011001111100001000100100010101100001111001001000110000000011101111000100110101111110110010101111001000001110110111001110111011110000010011100110111110000100110111001111001000101100000011000111011010010011011011011111000101101010111111110000011000001111000011110000100011110011001101101111110111001111000000010111011110110000011111010000001011000000000111111001000001110001000000111110000000000100100000000011110000000100101011000000011111000000000101100100000011110000010000001001010000001111011110000001000010100001111111111001111011000100000011111111010100000010000000000111111111001100000011100010011110101111011001010111000011111111111110010010010010110111111111101001110001101001001111101000110010001011001110000111111100100},
{784'b1011100110011100010111011000001100110100101101011110010010010111011001000111111111001011000101000100000010010000100000100001101100010111000100000000011101000010000011001101011110111011000111100011101001100010101111111101110100001010111011111110110111011001011111101101111011111100001011111111010011111111111111100111111101000111111111111111011110100000011110111010111111111100000000100011111000011111010100000011101111001100001000100000011101111010100100000100000001111001010000011010000000001110010101011111101110100000111010000001101101001110100101001001010010101011101111100000011000110000000101111100100100100101111000110011110100000001010100101010011110101010000000000010011101001111010010001000001010010011110111110111101000001001010101110111111010001100000101110010001000110000},
{784'b0101010110011110100101110011010010110100100010111110000000111010111011011100000110101101101000100000000100100001111111100000000000011111111110100100100000000000100111011001011100101101111011111010010100100010110011111101001000111101101011001111100101111110011111111001111011100001111011111100000011101010000111000111111000011111100000101010111111100011111111100011010011111100001111111100000000111111110001011111110000010110111010100000111111000101110011011000101011000000001101100001000010011011000000001111000000010000000000000111101100000000000000000000011001000000000000000000000111111111000000000000000000110111010100001000000000100111110010011101000000110001111011010000011111100001100111010100110111101011111111111101101110110111011111111111010111001011101111100011010011110101},
{784'b1110111011111111010110011111011010001110011011010101110111011001111111011111011001010101001001110111111110100110101100000100101111001011001110111000001111111111011011001110000100000000111101111001011101010100000000111101000101101000101000000000110000111100001000000000000000000000011000000011000001010000000111000001111000001011100000010010001011111000111101111111110011011010000001111111100000101111101110011101001111100011111111011101100111110101011001111111111110001000010100000001111111101110100000001010100111111111111001001110110010110101011111010000010111000000001111111110011000000100000010011111110001000100110001101001110111010000011100111110101011001100110011101101011011111110000000110110011100001000001000000000001100101001000000000000010100111001010110100000110000000010},
{784'b1111100101111011100101101110101100010101000111000001100010000100000000100110001001111010000000111000110000110010100011010101010010101000100000100010100000010101100011011111100100100000000100111000011111000000110010100111001010001111000111111111011010100110111111010111111101100111010111111011111111110010001100111011110010011001010011001101001100011000000101011001101001100000100010101001010111111110000000101001100111111111000000010001001001010100010110100101111110100001001000111101011010110110111110110111111001101110000111010101111001110010111101100101111110000011011110110010000101110011001101010001010001001101001111011110100110110110010011100011111110001011101101110010011100111111010111000010100011100100100100110010011000000000100000000100010111001110101000011111000111000011},
{784'b1101100010100110100000100100001000000001100010000100110000000001100010001010011010101010001100101001000000100001001000010111001000001111110010110001111111111111111000000000000111111110111111001010100001001011100011111101110010001000010100001111111111000000000010010000111111111110000010010110101011111111110111010100000001100000111111101001111101001110000000111010010001000000111000000011000010000111000011100000011110100010001100001100000011111111011001100100100000000111000011101111110010000101111110001001111111110000011111111001010011111110000111111111110000011111111100011111111100010101111111111000011111110110010111111111110000111111110110000111111100110010000100111011110011101111010000010000001110101110000011001000010101010100000000010001100001011110110000101001011100001010},
{784'b1100101000011110100000011001100101010101001000111110011111110010011111111110101110111101110111101001011111111110100110011100000011111010011111101000110011001010100100011101101101111111001011000000000100011011111111100000011111011110111111100000000100110101110111111010000000000001010111101101011000000000001000110100000000001000000011111110000000000000001000100110101110000000000010111101111011101100011101000111011111011110000001110000111101111110111001000100011001011111111111110100000001111100011110111001000000011110110100011101101100100001111100100000111110111110001111111100110010111011100000111111101100101110111010010100101010000010111100000011000000000000010011100011000000000000000101010001001010101000100101001011011010100111010011100110110001001101110111101110111011001100},
{784'b1111110001111011100011100101110101111100000010101101011111010010010000000010100111100110001000000000000000010011000000000111000000001000011001101000000000001000000001010111011101000000001100001001111010000000000011110111000101011011000000011111111110100100100010000011111111111110101010010000011111111111100100100001000011111011111111110100100000011111000000000100001101111011111001010000001111100011011111101100000001011110111011011110110000000011001111110000011011000100011101111111000011111001111000011111111111111110000110101110101101111111111000000001010101000111111111000010100100100000011101111000000000001011111111011110100000100100101011100100111000000011111101101110100000000000000010111110101000000110000001001101001101111011111110000000000100011010000101100011011101100110},
{784'b0011000101001010110110010101101110000110010110011100111100000111000101111011111111111111101100110101000001111010100101010110111111010111110111111100101001010000001101010000111001101000000011000101011111010111100110001110011101000101011101000011010110001101111110001101000111101100011111001110011000111010011011010001011110101010000001010110100111111001110001101010111011101010000110100000011111110010110000000101000001111101100110000011111011100000101111111100001110101110000110010111000000111111101000110010001110000011101011100001001010001000011111010000111001010000000001111101010001011011000010100111111110000101111100000000000110110000111111001100001000011011000011111110111101010011000100001010111111001111000001000000111010100110100000010011010100111110111110010010001111111011},
{784'b1110010000010000100110000100011111100001001100000001000001110010111000010010110001101001010000110001111111110000001101011011000011110111100010010000010000000111111111000101000101101000001111111111000000011111101000111111110001000101100111000011111111000000000011110000001111111101000100000000000000111111111100100000000010000111110110000001001100011000011111100010000011111111100001111110001100110111111100001110100011000011111111101100110101100000110011111010000111111111100000011101100000111111010111011000101111010001100000000001000001111100001011000100101100101110110001001010000100001000011001001101000011101000100011111111101111101011010100001111100001100100101100001011001111100011110000000110010010111010111110010010011100010001111111111011101000101110000000010101100010001010},
{784'b1001111111101010000101011100011000011001110100010000011010111110101010000010100110010101010110000011000010110110111111100010100000010101011111010011101110111111101111010011101110010011000100010000011111101110111001001011100101110111011110001000111010011100111000000000000011110011111001110010000000100110001001101110011000001100000100111110000011100100110011111000010000100111110000000101110101000111110110101101101100110100011001011111010001111111001100111001110111111000001001101001110101101110110100100010111111001100111100101101010100001010001101000110100100111010010000000101000000011101100001111000010110011011110100000100110101010111110111001110110111101101111110001000101101010000101110101111100010110000000000000001101000110101010110000010100111101110111110110000110110110101},
{784'b0000100010101001010100010100000110100011100001011110111111110101111000001100000001100000000011101110111010000100111100000011101110100100101010100111111111010011010010100100001111111111111001010010110000111111111110011100010010111111111111111111111110110101111111111111111111111100011111111111111010111111110001010010100100110011111110001101110100000000000111111001100100000000000000011001100001001000000000010001100010000011010000000001000110001001100011000000000001100000000000001110000000111110001111010100011000000001110001110000110011111000001111111110101000001111111001110111111000010001111111111001111111100100000000111111111111100101101010000111111111111100010100011001101101111101100000000010000001100111111011110110100111010011010101111010000010010000000111000000000100000101},
{784'b0110100010110110011111010111110101011000101011011010101110100001110001100001001001111100110010000000000110000011101101100000000000001000001010111100011111000000000011111011101000010111110101100011111110010111110111110010001101000101001011111111111100101110100101011101111111110000011001111101111111101010101010110010111101011110001011111011111111000100101100101100110111111010000000100110010100000111011100000111111101101111111111111000011100100101011001011100000000000101100100100101110011001100010100100110100101011100101000100011101110000000000000001000110010110010000000000000101001111111110000000000000100001010111010010000011001011011111001001000001101101100100100111001010100001101101111110001001010011011000011110111010110000111101111010001011101110101110111111111100011111010},
{784'b1011110110000101001011011110111110001111010001111011101111111000001111110101101111110110011101111101111001111111101011101111110100000001110010000100100001111000000101010110101000111111100000010101010110000001111110000000111111001000001111111100000001000000101011111100111100000011111010111110001111111000000101000111110001111111101101101001011011000111010100000000111010011000011111100000001110000001100001001100000001101111000010000101111000000001000010000111010010000000100101001000001011000000000011101111010000110000001001000010110000110110100010111111100111011000111100001011111110001001111010000011111011111001111101000011111101111111101111000000011011111011111111001111110001111111110110111100111010001101001111111111001110010011111111101111011011000000111110010011100100110110},
{784'b1001111111100011110011010100011010010001111010001101011010100000111000001101100011100111110000000001010000111010011101000110111111111111110011000110111111111111011101100100010100111111011111011010000010000010010011111111111110100111111000011110101111011101011110000001110101011110000001000100011111101111101001111111111111111100000010000110011111111110010101000011100111111111100101001000000101101101110110110110000010100010100000000000000000100011110100000000000110000000001100011000000000000000000110011111000000000100000001000001111000000001110000000101011000110001111111000000001010000000111111111101011011100100101101111111111111101101010100101111111111111111110000000110010111010001111101111000101000000000010000000101000010100001110000011000010110101000010000001100100111001010},
{784'b1101111111111010101001001001111101001000010000100001110101111111100000011101010111010110010000000000000000010001111001000000001100011101001100000111101011110000010000110001000100100111111101000000100100110111111111001111000111000010111111110101001110101010010111111000000000000010000001011001000000110000000111100011111100000111100001010011111000000001111111110010000111100001111111111100010111001111101111111101000011111101101110111111110000110101101001111111110111000010000111100011111111110000110110100000001101111100000101000111011010001100000000001110010110100000000000000011110100101100000100000000001111111100011001000000000000111100010010000000000000001111001110100011000000010011111111100100001101000001111111111100101001111101101010111110101110011110101111001110111010000110},
{784'b1110100111001000011011001101101111001111001000011001000100110010100001101000111011000011000010000001011101111100001000011110110001011110000011111111101110110100001010001011000010111111110010100011011100101111101100001001100010011101000100000001000010101010110110100000011001010001101001101100000000010001000011110111111111000100101010101111101111111000111001111001110111111111110011010111100100011111111100001001111110010010101011110000010111100100001101111111000001111110010011110011111100011111101000001100011100100000111000000101000000010100000011101011100011101001010001001110010011000000000010010001000000011011000101111011110100000001011110000010100000000100101110000110011100110000000110110001100110011111100110111110011110101010111000100100111111011000100111011100101001011111},
{784'b1010110100110011111011110000011010111011101111101011111100101101011000101011110001010100111100010100000001110011010000011101100111001111000011110001110000100000000010111111101101001000000000000111010110011101000000000000000111011011001000001100110000101100000111100000001110100011010001111010000011100001110111001010011000000001001111110001110110100000001011011101010101011111000010010101011110110111100111001111110010000110011100011111110110101110011001110001111110000011111111110110000111111110000010110001001100011111110000111101000001100001111111101111111101011000011111101110101111101101010111111101010000010100010100000010011010111110101011111010000000001111111111111100100000001001100010010101010100000000000000110011111011100110001000010010110011101011010010111110100111001001},
{784'b0000110101000100001100110001001101001101110000011011011000100000001011101111000011010011100000111000010000000010011110111001011001000111100010011101001111111000000000001100001101111111111100001100101110101101010111000111101101001100001000111010111110111000011110100111000110100100001111101110011101110011001100001111111111110000111110001100001111111111011001111000011101111001001011110011101100101011111101001011110111001011011000011000011110100010011111111011000000110011000011000100110000001111111000111111011110010100011110100001010100110010100011000000111111001110110001100110001010101110101100000000000000001001000010000100100000000001110011100101101111010000011000000010111100101110010000110111001001111111101100011010100011011110110101111111111111000101000000100100110010100100},
{784'b1000010000110011011100110100111110010010011001101001100001111011101011100100011011101001101110110100100110101000000110110110001010011011110111011110111101110100011111000101001011111010000010011010000010111111100001011101111111101111110110000000110011001000111111110000111110100010101001001001000000011110001100001001011001011111110010010111011111111000111101111000110111111001000111100111101101111111010000011100011000000011001111100011111111110111101000111100000110000011100101000101000000111101001000111000000000000100000001000111010111010000000100011000011100010110100010010010100010001000011011110110011011001110111101111111001111111101011010110011001101011100101001011101101111010000100010010001100001011110100001000000000000100111001000000110001111001111000011000111011111011010},
{784'b1011111001010000100100001000001101010010001011011011010001000100101100000101110110001111010101100110111010010011001100110000111111101111100111101001000100111100100001100111001100110010011101100111000010000101000011011110001001100011111000000111110011100111001111100000100010010111101010111111100011011111111110111011101110100111110000101111101100111011100000100110000111110101110001100100111110111110000111110010101010001110111110011000110101110001000111011010000001001111001101111100000000110100010000110001101110100000101001101011011001100000000001111110010011011000000000000101001000011111100001000100110100001110010110001000000000101000100110010011111000110101100000100100111011011110110100100111001111101111100011010011101000111100100001111011000100010111101001001010001010000111},
{784'b0111000010000100000011100000000001000101001010111110011010011010110101011000011111101000001101101111111100100010010101111011110110101001001100110100011100000100011000011010010010100000011101101011001000011000000011101110110101000011011000100000010001010111100000101111000000101100100100111111111100000101010100111110000000000001100000001011000000000000101000001001000000000001011111111101010111010000000001111001110100000110001100010111100100001111100000010000011101010101111111111100000001111000010111001001110000001000000000011100011100000011110111010101111101101100111111000000111111111110000111110110101100110110000101111111100000000111000101100111111000001001001011000010100100010110011010110100100110100001100101100111001001000010001001101100101001111010010101011001001100100011},
{784'b1001010010110110110111010000111111001111110001001101101100111000011010000100110111011010000000110001011101101011010000101000000110011101000110111100001000010001000110111100110111000001010101101010101100110010011111000110100010001111110100110001000101001100101000001100000010101010000111011100011000011011000111010000101111111100111100011111011111011100111011111111001111110101000111101111000110100011101100010111111010000001101111110000010000110010010000111011000001111101010100000001111110000000010100011000011101011001111001000011000101011011100010100000000100110000010011110000100000100101000000000100010100000100101010011001111110000000001001011011100000000100000000101011101011011101110010001011110110110011111111011111101110001110101111101011001111100010010111101000111111111111},
{784'b1010001010111111110011110011101110011010001000010010101011001001010010010101101101100110000100111000011001001111001101110000000111101011010111100110011111000010101100001000101110111100001111000110111011100001110000111111001101010011011111000011110111000111001001111100011111010011100100000001110001110000101011110110000111000111100011010101000101111100011000001100010100001111100001110001111011101001101000001110010110100110110001000000000101010101110101111000000000111111011111000110010000001011100000100111111100000000111111101001011001111100011001010100000011101111111111101011010001111100111111111110010011101000001100010111011111110011011000110001101111110000000001110010110100100110000000101101111011000000100001001011110100101110010000010000101101000111111101111101001110111111},
{784'b1110111111011011011110001011010010110001011101100100111110110111101101111111011111100101010110111010101011110101111011000000001001011111000011100100000000100101100110011111010000000000000001110001100101000010010000000101110010110001100101000010001101011010000001001000000001000101111000000001100011111101001111011010111110001110010101101010111111111100101101001001110001111111100001111101101111110111111110000000111110000100001111111100000100011001100011111111100000010001000001110101111111011101000000111111010111111011111000000110110110100011001011100001101001100101000011110000000001111101010000010111100000010110111101000000111011110110000101110010100101110010100000111100000101011101100101111101000110001001001100101100110110011100110110001011011010011111100101001010100101100010},
{784'b0010100000110111010111101001000000001101000111110000010100100111100100100010011110000000000001111110010110011101100001010110111000110100000111111000111000000100000000000111010011100000110101000001000011110101110000100100000110011010000110001000111100000000111001001111111111011111000101100111010011111111000000111101101000000111111110000100101111010000101110110011000111010010000000000001100011101111110100001000011111100011110111110000000011100010110011111111100011111011001110101101111101011111111011100001000011111001101100000001111010011011110001000100011011000010001011000000000010110000011000011100000000011101100101100000110000000001010011000001100000101100000011010010001000000111000001010000100101111001111101110111110010010011011111011100010000111010001000000101100100101010},
{784'b1111100101100111111101110111100000100010010001011101110110100111101000011000010111111011100100100001001010101111011100100111111101011000001010010010001001011001101000111001011110011011001000001001111001010100101100000000000010111100111000000000000000110000001100000000000000000001011100000000000000010000011001001000010000011111000011111111011000111111100000000011101000100111111110110000101110011111111111111010101111101101101111011110100001000111001111110001010110110101100111011000101001100011111010001111101100000111111111101001011010000010000110111111111110001110000001001111101111111011000010101001011001111010100011000010110000100111010111010100101000100101011100111110100001000111001111111101101000100000010000001111111110101111011001001000110100001100101011100101111000011000},
{784'b1111111101100100101111110001000110001100100010001000001011111111110001101101110011101010010111100000000000011011111100001110011110110111101111010111111000000100001110001101111111000000000000011101110111111000000000000000110100111111110000000000000111001111111011010001111111111000011011111111110111111111100011000110011110011111111010100110110111111000111111100110001011111111000001111111111111101111111100001101111111001010111111110001011001111001000101111100001111110111001100101111100000111110011111101000010000000011111111001001110111100000001111100000010110000001000000110000000000110011000111000100101000000011110100010100100101010000111001010010110011111110110001010111110001000000111101011110110001100000000110000000111100100010000000010001001111101101100000000011100011110011},
{784'b0100111011101000111110011100111101010101101011111100101010111101111111011011111100000110100010111101011111001111010111010110111111010111000101100111000010001100000001010110110111000100001000101011000010011110000011000100100111111011111111100000000000110111110101011110000010001010101110001110111111001001100010101001000111111111010011111101010100111111111000000011001000001000000110100001110110010000010000111000100110010110000000000111010011010010000001011100011100110011000011100111000101101010100010111100101011111111000111001001011001010111110000011000001111001100000111100001000000110000100010111110001110000011010100000000011010100010000001010110000001110110000011010001110011100111110100100100001001110111101101111101110000110000011101111011101001110001000000011101000101110011},
{784'b1101110111101001000000111110011111110101010111011101110110100000010000000101111111111011100010100000100000011101100101000000000000010110011011100100100000000000000111000100011100100000000011111101010011011110000001001011011110011100000010001010101101101111111101011101111111011010010010100000001111111100010101111011010011011111101001111111101011100001110000000101001110111100000101001110100100111111111000001011000001110111011111100011100010011011111110010100000111100000010111110110111001110100100100011110101001001111000100010111011000010001101100000001011111100000000000000000000001010110010000000001000010001011000001100101000000001110110101110010110110101010110011111111111001000001110011001001111011111001010100000011100101011100101101100001001110110101011001001101101110010011},
{784'b1001111100101101001010000110000101110010000011000000000010100011100111000010110011001011000111111111011101000000000001011111111110111000000101001111111101111111110000000110111111010101111101000011000001111101101000000010000011010110000010000000010000110101111100000011001001100001000001110000001100001000010100101010000000110011010000010000001010000011010000001000100001110000001111100000110101010001010001101010000001000010001111000111101101110000101101100101110111111110110111110100001111000111111100111111100000111110101101110111100110000111100011011111100110011001010011111101111101001001101110111101111111110110111101110000000111111111111000011111100000011110010000001110010101001111001000010110010100111100100010101100100001110001111011011101010011000000100111000010000010010011},
{784'b1010100110011001000100101101111110100100010010101111000001000001000111010000000011000000001010001110111001100110011100000011111110001101001001011011011111111011101101001101110011100110101111111101001101110110000111100101111100100000011010100110011111010100100011111001111011100111010110001111110010011010111100110010001111011111010001001101000001111110111100000011101000000001111011010000010111011101110011010110000000000101011111111001100101001100010111111111100000001111110001011111111000000011011100001010111111000000000011111010000111111100000010010111001001111111110000010010111100000010111110000001101111110100010101010111100010011011000010010111100000000000010011000010101100110100001000001100000000101010000000000101000101101011001100101100011001010110110100010101010000000000},
{784'b1011101000110011001110001100110100011001100010001001101001100001000001010000110011000100001001101110110100000101001111100111100001110101001011100000111011000010100001101111100011100000001000001011110100011100010110000001010110100100100000110000000011001100011101000011000000010011100000111100000000111100101100000111111000000001011000010001111111100000001111111100100011111111100110000111111111000111111111110111111011000111010101111111011011000111100110001111111111100100111111001111111111111111110111000111011111111111111011111111010011011101111110010111101000011111100000111001010101110011100101000111000001110011100100001011100100001111101100010100000000000010111110011000000010111100000110011100110110010000001101101111101111010110011010111001010100001001110111011101010000001111},
{784'b1110111101111111110111111001111111111100111100101101111001111001010000010110110100100101011110000100000001000001111100100110000010110100101101111100000000100100010111101110000000000000011111010111010000000000000110111111001110000000000011101011011110110111100000011111100111111101010010000011111110001001110100110000011111111010100011010101111101111111010100111101100110001000001111000000011111110100000001111000000011000111100010000111000000000110101010110111011100000010010011111111111111000000000001001010000000111100000000001011111100011101110000000100011101000000110110000100010010010100101000001001010010101111011100101001011101110000111011010101000011111111011110011000110100000000001101011110110110010110101111011111101011100001111111111101111110100010100111110111100110111101},
{784'b0100001110100000111001001000100010000011110100110001000001110000110110010011111000000000000010100111010111000000001001111101010111111110110000111110101001100100011000010011010111111011001101111110010101011111111110101011110001011011001100110011011111001010011111010000101001111100011111111010000011110111110001010010110111110111100010100011111000111111001110000001010101001011110010010010001100000010000011001101000000110000100000000101111001110001101011000000001101001001100011001000000011101111100010001110111000000111000101100000011101000000111101010101001100001010100111101111011110001000000000001001110001001000110010001000101101010000000100000101000111110001011010100010001101001111111011001001101010111111111111110000101100011001111000110010100000011010000011000010101111011111},
{784'b1001101100000100010101001011001100000101100101010001000110000101100000011110010100000010010001010001100010101010000110000111101111100011000101000000001111111111110111000100010110010111010111110100011000101000111001000001110000001010110101000000000111000101011101111000000000111000010000100111100000000000100010000011111110000010000000100101001111110000000110101100101110111111111111110110110000111011101111110010110110111000111101110111100110001111111001001111111111011111101000011110011111100100011010010010011111110101101101101101111001111111110111111111111001111111111111011111111110000000011101111100011111110000000010001011011001111111010000011000010110101111111110000001010010111001100100010011011110000000000000000010001010000110001101110100100110101011100101110100010011001010},
{784'b1011010011010111011011010011110000110100011100101010111010000101001010100011110000010110010001000000101111101111011111010111001000000000011011000000010111100000101011100000000010011111000001111100000000111000111100001111111101100111100111110001111111100010001111111110000111111111110011111111111000011111111011011111100111000011111011000101111100000000011111000110000011000000111101111100001010000000000111110011000000001100000000100100001000001100010010000011100011000010010011000000100111100110010010000011100000111010000111000101001101000001111010000011110110011111000001101010000001000111101011000101100000011010000000100100101110101011001000100010001100101001111100011110001000000010000111100010111100101101100110111110111000000001011111111111101101100110111110110111000011001101},
{784'b1000000100100010000100110111110011001101010100001100010110011101101111111001011011001010010110101111111000101011011001110011111111111101000011110000010010111111110010100100110001000001111110000100011000000100001111110100110000110110110110011110010000110000011011101000111100001010101001111100000111110000001001011111011000101111100011010010011000000011111101011010011100000000010111111011101000110000000000011111000111011001000000000010011010000100000000000000000111110000101010010111001000000000100100110000111111111111111100001100010011111111111111111110000110001111111111111101000010000100111111111000010010100000100111111101001111111000001000101000000000001111111100010010000000000101011101111110110100000001000101111100010000000000111111111110101001110001001001100000111000000000},
{784'b1110000110100100111010110110111000000010000000001111101000000000100000011000110001100101100001110011010110010010100101010011100010110100010001010011111100011111101110001010110001000100101101111011001101100010101010000011110011100100001111111000101110101011111110100101001000111000100011100101110000000101111000000000001010001010000111001001000100111000000000000011111010111110000001101000000000011101111000001000110011111110111111001000000010011000111011011000000001111111001000111011100000011111111110010111111101100001111111100110111000111001001101011100011011011110101101101111011101010010111001111011100101111100010000000101011111110101101101100000001010010110101011100011011011001111011000110101000100000010000111100000000000010000111001011101001000010010101011000110010010010110},
{784'b1111111101111010101111111001100101101111101100010111000011100011111100110111101011010011001010100011111111011001001111110100010111011111101111001110000000111011101110111010011000001011111111000011100000000000011111110000111111100100001111100100000011010100101001110100000000000010111100100111100000000000010001101000001111000000111000101110101001110110011011100011011010000100000110011011110100110110000000111000110001111101111000000011111110000111001001011100111110010110101000000101110101111100010001100101000101111111110010110010010010000101111101010101100100110100010101011001111000110011110000100111111110001000000110010100001010001100111101011011001011010011000110101100101101111001110011011100001000101011101111011111111000010111110111111001111011111110111001111000111111011100},
{784'b1100111110110110000000100000000111001101000011000000000110110111100001100000011110001101011110011011011010000001001011001111001100111101101111100011111111111111111101010010110001011111101100101001111010000001111111000000011100000000000001001000000001100001000000000000000000000011110000000000000000000011101000000100000000111101111110001000011110011111110111111101000011001111111111111111011100101111111111111110111010001101111111111111110110001100001111101111111010000000100011011100111110000000010000101000011111100000101101111001100110111111100011101111011010011111111100101111111110001000111111110010011011110010001011001001010001011110010000011000110110000010101000000011000001100110100011110010110000100000001000001000010000000110100000100100100010010100110101011000111001000100},
{784'b0100010101000011100010110011100001011111000011010010111001011010000111101110001011001010110010110111001010111010010100000010001001011111000000111010100111111111000011011110001100011011010001011100001110101011111101000111001100000000111110000100000001001011111011110100000101000011001101111111100111111000100100001111111000000101010111001111011001000011001111101111100111111101010000111110111100110000001101101011000011001100100101111111100000000111101100101111111111000001111011100100111111110000000011101010001011111111000011111110001100111011111010100011101100101001100010001111111110110000111101100011010011111100110000101010110000111111111010101001100010101011111000000011100001101110101101000100111100010000001101100010011010101011110010010110101111101011001010011100101011001010},
{784'b0010110101011001001100111000001001000010001110011001011110111001100111101010000001111110110010000000101100101010101111101101001111111110101000010111110100110001000110000010001111100101100000000011110111111100110000100000000011111100100111000100000000000000011110001111111110110000011111100000111111111111001010110111000011111111111110111011100000000001101111111011100110000000001100001111101010000110000001100011101011001101011010000011000011100000001001111100000100011011000001001011111000010001111100100011001111111111101000000101111110110011101001000000000011100000001100101011010001011001101011010010101000000001110100000000001111011000010000000011001011000111000001100110111001100000000100100111111111100000000100000000110100101001000000000100110101010011001011001111101101110110},
{784'b0010101111010001001100001100111000101010100010011100011110111100010011000011001100110010000101101111101000010000110011011001100010010001000100111010000000000000000000111100110101000001010000010101010001010000001000001010001010111000000011100000010001011111010000101111111010100010010111010000011110000000001110111000000000110011000100000001000000000001101000010110111000001100000011100001100000100001111100011100000101000110110110010111111101011001111101110111011011110101111111011000111111111111101100100101110101101111111111111110011110001011111111101110111110011111100111110001100011101101101101001010110100001000010100011111010101001001110011001111010000010010000101110111110111011000000011000111000110000111011000010100100001111011010000101010001001011000010001110111001010111110},
{784'b1110010000010001100110000010110001111101100001110010101001000001111110000011110110101010100100000000000101010101010110110011000000010100110101101100010100000001111111101100100101000000000100111001010000100000010000000111111001011000101111100000011111001010111111111111000000101100000001111111111100000001111001111111111111111000000011011001111111111111110000101110101011110100011111100111100110110100000001111100001111000010000001011111001111111100101101101000011110001011101011111001110111100011111110001100001101010010000101010000001001101000000100100001001001100011100001111000000000000100000110000111010010000000010010100000101101111001001000100100000001111111100001111111110110000011101100011110110101011011000011111100100110101111001100110001110010100001000001001100011100001100},
{784'b0111001000110010000101001000010010010000000000111000011010011001001101110000001101001011101111111001101110011011010111110001111011011010001001101001011111011111110010100100110001001111111101111100001100000101100100111011111000110110101111111101111110100011000111111111111111101100100000111111111111010111000010101111111010111111011100101001101111100001111111110000010010001100001111111111100000000100000000011111110110000000010101110111111110000110001000010101011110111100101000000111111101111111100010000010111000001111111110001100000011111111111111110000111010000111111111111110110001011101100111111101110110110100100000001011111111000111001001100001001011111011011000110000100010001110101000000110000010001100100001110000000110001100111001011101000000001011011001010110100100000110},
{784'b0100111110011101101111101111110101001111011001001111100110111100001101111001001010110111011011010000100010011101110010110111101010001001100111101101111111111000001110111001110000010000000011110010011100100000000000000011000011110100000000000000101001111111100000000000100001000010010010000000000111110100001101100000000000111001001100110111000010011111100111101100001001101011111110101111111001010110011111111111011111100011111111111111111111111110010111111110111111111111101111111111110001111111111111100111111111000111111111011101011101111100001111100000001001010101100001001000000000001101100000000010000000001001101101000010000100010100011011111000000000000000110001011101101000000000000000000011111111000000000000000011011111010100000000000000001000111011111001111101100111101111},
{784'b1011001000000101000001000010010000001100000100000000110000101100010010011000000000000101000000000000001110110001000111100000100000111001101101010011101000001111111011100001101000000000111110111000010000000000000000100111101100001010010000000010110011110100001100011110000011011101000001011111111100011011011111101100111111110001110111101011011111111111000100110100101111111111111100110110010110001111111100111100001000000001111111000110101111111100010101111000001111111111011001100111000000111111111100101010011100000011111111000010110011111000000111100101100011101111100000001111110101111111001111100000110111100010000100110111000111000001000001100010110100000110110100101001100001111001111110000010010001000101110001111100110010010010000111101110100101110101001001111001001110000000},
{784'b1100011100010110110010110101111011101110011111001001010111001111011110111100011111111011101010000001111010001011110100110000101110000011010111010000001011111111101100111110000001001111110011101001111110001011111000001111011101000000101110100000000010101010000000111001000100010110011110101111111100000101011101110011110001111011100011111010011111000011111101110011101111111100011000011100001110011111111100000000000001111110100011101000000000011011100001101101000100000000111110110001111000100000101001011110110111100011000000101010011010001100010010111100111101000100110000100111111011010100001110101100101011101110110010010000101011101101100111000110000010001000011100001100001000000000011111110111111101010000000001111110001011000101111111101011101111111101010101011001010111100010},
{784'b1100000100000001001100100101001101110111101101001111100000010101001011101101011011000110110101001001111011111110101111101010111110111000111101110011100010110001010001000010101100000000000001000010101111010001000000000011101011011001000000000000111101000010000001100001000101111001001101000000011111101111000101001000000111111100111100010010010000001111111100101100000011000011110010111000110000100010011000111111100000110111011101001111111110100101011100111001001111101111101100001111111001111111011001100111011111111111100000010101111001111111111101000001100101001010111101110100010001000001100011110000001000010100111011000011010000111110110110010100000000000111101011010100100100000001010001010011110111000000000100000101101100100101001000001000000101110110011000100111111110011111},
{784'b0011111011000010001011000111011111000000000001011010010000100110001000011110000110111110000111101100000100100010001001110000000000010011000010111011110100000000010111111110010000111111000000011110001000101111111110000000110011000101111111100000000011001110111111111000010000000110001011111111000001110000011010001110100011001101000000100111001000001100000010000001011010010001110000011100011110000101101011000100001011100010100000101111111101111110010000000001111101111100110111110010000111111110111000011000110000011111100111100101110100000001111100110101011010101100000111111011111001110011110010001001111111111010110110010000000001111110110011010111000000000111111011111101001101001010100101010111101000110000001101010111100111111010000000001001010101101101000001000000011000011001},
{784'b0100101100001000001101000001000000100110101011100100110111110000101001000001000110010000110011100010111011100000110101111011100100110111110101111101110010111100110101011100110011011100011111100100010011110101111010011110110011101111000000011111111000110000110110001101101111110000011000000000011111101100011001111001000001111100101001000010100001011111110010000011010100010000111111111100101101110000101011111111010010010000100001011111111110101100011100100110000001111010000111101101111001101111011010010001101111100010110111000011110101101100011110001000110001011101111000101000100001001110110110011100000010100001111010011001011111011100100001111111101111010011100110010011110111110101010001110011010010111111111000000011010000110110010111000100110001101011010010011101110110010000},
{784'b0101100000000100001001010000000100101011101011101011011001010110100110011000001001010011010111110101100001011000001110111111111010001011001011100101110110110001000110111110101111011000000000010011011101111111000001000000000001111111111011111011000000011111111101011111110111100000010011111111111111111101000001100011111111110111111100001011010111110001111111111011111100101000011111111111110100111001100001011111110110011110001011000111111111100100001110011111111101111111110100010000101111101111111111111010010001111101101110101010100000000111100111101101100001100000010010111111010000010100000000001111111101100000010010000010001001100100111000100110100010100010000101000111001110010010100011111101111010101111101000110010001100000101000000000011000001100100100100011010000001100010},
{784'b1110101111100101001000011111100100101110101101111001000101111110101111110011010101101011001011110001110100100010010000010000000010101110001011101010100001101011101011010010110010110010011101111101101100000010011000000100000010110001001100001101000110100100101011100111111101000111111001111110110110111001101010100011100001110100111001110101111100000011000011111011010011111000001000011111110100011111110000100000111101010100111111100000000011111000100011111110001000001001101100000111111000100001111011111111010111100110001110100010110101011111101001110010100011010011011100101100010101010110010011111010101111100101010101101100111000100011000111100111010010001110101101010000010010000100101000110101101000100000010000111111110010100011100011101111101000101100000110110000011101000010},
{784'b0100001101001101000001010101001000100000110000011011110011011111000101010100100000001111001000000111001101001110001110001110110100001110111000110011011000111111111100111110100001111000001101110000011100111001000000010111111001110100101010000001010111000010111001111100001000011100101001100111110011011100011010100110101000001111000100000111000010100000000010001011000000010000000001011101101000000000000000100101100010100010000001100110110001111111010010100000101111000111111100100110110111100110001110100100111001011111000100111110000111001111111110101111110011101100110111000101011101100001001110000011000011111010011011110111000000111100110010110111111010101101010011110000010000100111111000101101101010000000010100010010111111001001100100000011010111001101110111011101011100110110},
{784'b0000011000011101011011101011010111101110111011101010011010111000001001010000111111001011101110001000000010001100110010011001100010100101101100100101001010111111111001101011001110011010011101110001011010110000000101111100110111101011000001110110101101010010110001000111111111110011011100011001110111001110000100101000001111110010101000010111110110111000111101110101111110001111100011001010110100000101100100000001001011001101100001000000001110101111101010010100000111011111101110001100110000000001111010100011111011000000000101111111110010010110101010000000110001010000001010000100111001110110101000000000000110111010001000000101111000011001100011101011010100010111010101000111111010101111101000100001100110100000101010010001110001111100000000001111100110001101000110100110100010101010},
{784'b0010000100010101101101110011000000010100111111100100111000011101000001110111110000110110110001100000000000110101100010110000000000000110000001010100001000000000000101101111000100100010110111001011100100010101011001110101100001101010001110011110011100100010001111111000000111101011100100111110010000000111110001111111110001000000011111110101111111000000000111111111010011110011000001111111100100010111111110000111111111100001111111101001111111111000100101111011110111111111011011011101011111011111110110011110000011111110110100001011100010111011111000000001011100000001010010001100000001000100000001100110000000010010010000001100000100000011000010110101011000101000001101100101011000011000100000100110111001100011010000100100101111110110000011010101001111101001010101000001010000110001},
{784'b1110101100010111011111101010111000110111010110011111011011110111100100110111111101111101101101100000000001110011100011110010100000010110101111101000000111000100100111110111010110111110001100110110001000010111100001011011110111001000101111000111011110011111000001110000110111110100111110000100110011011111010100111000000011111100010000000111001010111111111011000011001110000001111111111100010101001100000111111101000001110110000000011111001101010001101010000000011011000000001111100000000000001101000000001010100000000001011000000001111101000000000010110000001101111010111000001111000010111011001111110000110000000010010110111110000101100000001100111111010000110000000111110001111111100001100011100011111111111110100000100011101111111111001000110001101111110010111100010111011001010110},
{784'b1111011011011001110100101110011011100010100011101100101011110000010110000010111111111000110101111110110110010101101011110111100000011101111111011100011111010100001011011011101111111110100101000011001000111111111100011110100101111111101110111100011000100001011111000000100011100010001100000000000011100001001111101000000000000010010010111101000000000000000010101101000100000000000000001101100101010000000000000000111010110010100000110000000000001110110000001111111000000010111110111011111111000000001001101001010111111100011011011100111010111111111001001010010101011111110111111111011100100101110111111111111100111011010111101101001111111011111011111111000101110001111001000001010010000000111011011100111000000000010100101010001000110100011101110100011011111110010010011011110111000011},
{784'b1110000000000100001100110110001101011000000101111101100100101111010010100001001100000000000000000010000101000111111000000000000001011100101010101000010001001010111000000111110111111100011111101000001100001101110111011001110001000110111000110111110111101111011100001111000010111111001101001110111110001011110110100010110111111000001011100110111111001101000000100100001001010000000000011110001101101000001000010001111111001101111000000000011111111000110010000000000000101111111111101110000000000111001000011101011000000011011001000111111011000000100100010000000110000001000011101000000011111110110110111111000000001000001010010111001000000001101111100111001001011101001110010011010101010001011101010011000110011101111101110100101110001110100000111111100100101011111110100100110111000111},
{784'b0001011101000101010011010110100100010000111010000100000001000101000101001110000000011010101100010000010110100000100101010101101111111100010010000000100000111111111101001000011110110000001110111110010011111101000000111110101111001001011111000011111111000000100111011100000111111111110001011111100000011111111000100001010000000000111111100001001101001100000000001110000000010001100000000001001101100100000000100000101110010010000111000110000001011100001001110100110000001111111111011111110001000011111110111110111110001110011111111100111111111111111111101001011110001111111111110011101100010010111111110011011011110001010011111010000010111111001011100100011011111111111000001100101001111111000100001100011000000001110110000000000000101000000000000000001010110101101010100100100100011000},
{784'b0111000010011000111111100010111001100010111001111001011101000111110111000010110110011010111000100011110010000101101110011111101110100001111011111111000001011111000000110110100100000111100010100001000010110010100100111010001001100101101100111111101000010010011110100011111101100000010111101000001111101001010011001000000001100111101110001111000010001101001001001111001100110000111010110101111111011110010111010101011101011010101101011111100110110101010111010001110001101011100111011110011010000101101011110111100100101101110111011001111010010011100111101100110011111101011000101111010000101110100100101001100010010111001011101111110100000001011111100001111110001011001011111010100110101111001101101001110110100010010010010000101100010101011100010111101010010001101111100111101111011110},
{784'b1000101100100000001111100110010001100100011100001101000010010110100001001001011100001010000111111111110000101110100001011111100111000100010011101100111111010010010000110001011111111010111010000100000010111100000000001010001010001111101010001111110111001001111111100001111111111100000011111000000111111111001000010111110100111111111110100100101111000000011111111000001000110110001000101111101100100001000101100000011110110000001111011110010000001011011111001101110001000111110110000100100111010001011111010001010100110000000000001101100001000111000000001111000011000100111111011000011100010000000110010100000111111000101011111000000000000110010001000011111000010110011100110000100011000010111110000000000010111110001001101010000001001110011011110111110000010111100110010010111010100000},
{784'b0111110111011001110111100001010011111001110011110111111101011111000011000010111101100101011001111011100001001010101000011111010100001110111011011010000111111111011110100111111000111111111100001001011010000101111111011010011110001000010000001010110000001110010100000000001011101111101111101000000111111111111010000010100000000111110011001001000000000001100010000010000011000101100001001000011100000000000110010010010000010110000010110100000100101100111011000000011000011001110111111110000001011100000001011110101010100111111100000110110101100101011010011010101000001111111111100110001010000111111111101001000000100000111111011111001110011111101111011101011111001111111111001111100110001111111011101101110111110100111000111010010010111001101000001001001001001111011101110100011111010011},
{784'b1000001001000010000101000010111001110010110011101001101101110110011000111010011111111001110010001001010101011100010001010000000001001110100101001101100010000001001101011000110011110000000000001011010101111111110000000000000011011111111111100000000010110101111111111111000000001100010010111111111110000000100100111011111011111100000011001000011100011111111000000100101010001011111111110001100101010000111111111100011101011010000000111111100101111111111000100011111110011111111111110001000111110000111111010001010000010110001111111100111000100000000000000111000110011100001001100000011000011110111000011000000010000001001110100010000000000000011010000101100000000000000101101100000111101110000001111010011010011111110100100110100010100010110101010100101100011101110001001001010011000101},
{784'b0011011010111011100111010101000110111101001111101110111011011110101100101011111010111111010011000000000101001011101100001011101000010001010000010000011010110001111101101110110011011010000010101011111001000010001111111110100101100001110000011111111111100000101010100000100111011101100010101110000000000000011011111011111100010000000011111111001111110001100000000010110111111111100111110000000111011111111110001111100000111001011111111000111000100100010001001111110100110100000001110100111111101101101010011100011001111110000100001010011001010101111101111101111000000000000011111110101110111011000010000001011111100011111100000000000111111111001100111000001010111111111000100011101001010001011101110101110110100000011100011011000010000111101111000111011000011110001100100100100010010001},
{784'b1010000100110010011100011000001110001101110011110010000000110101110101001100110101001110101011101111110110101000111011011111111111110010010101100111000011111111100001111010011000000111111010000100010101100000111111111100001101001000000000111111111000101001000100100011111111110000000001000001000000111111000100000000111000001111111110101110000011100111111011111000111101000110111000000000011000000110110011110000000000010111111000011110100000001110010010000111100010000000001001111001111000001000000011101011000111100000000000111110101001111110000001110101100110001101011000111110010011100111111000001111111110011001110000100011111111110001100110001101111111111110111011110010011111111111110000000110101110101101011110101110001001010010111111111111100110011111101000100111000001011111},
{784'b0011001111100111111001011001001101111001010100010101110111111110110100101010110000011110001111000001001100011000111111000001100000010111111101001001011111011010001000111100110010101010110100111101011011011111100000110011101001111110111100001100110111101101000001111000011100011100001010111111100000111110101011101101111110000110110010111011011111111000011011100010010101000111000001001010101110100101110100000000100000100111100000001000001011000100010010000000100001011110111111001100000110000111101000110110000000111000101101111011110011000011100001000010111000000000011110000001000100110000100001111101101001001001111010101111101001100110010001111110001110101100000101110101110011101100000010111111101001110000100110110100011100011001010110011000111101110111101110101100111011100001},
{784'b0010110111110000010000000110101110110010100110101010101101101010101100110011011001111110111010010010001010101110100110011100110000000111111100111011111111000000011100110001110111111100000110100011100000001111100000001000000101101001111111000010011000100011100101111110011110000010010011111111110011111111000010111011111110001111111011110111110111110000111111100000011010010000000011111111011100111110000000011110111101000100011000010001011110111110010010010000101101101111111110100000000011110001100011011101000000011110000000000100010000000001111000010000010011000000000111110001000100001110000001011110100000011110000010001011011110100000100111000000000000010110001100000001110000000111010100010001011011111000010111111010001000101001111101111110110110010101111101001110000110010100},
{784'b0011001010010100010101100100001000110001100010011101111100000000111010110010001000001000110110011111111110001100110011011011111111001101001110100110001010101011000000000010110111000101011001111100010110000010110110000010100011100000010110100000000100110111101011111111010111111010110101001011111111111110001001111110001000000111111110000001100000000000011011101100011010000000000011110111101100010001000000000001000011000110001111000000110110000110010011111000000000010000110111101111111100000101110111111010111111111111111100101000101000011111111111111011011011100011111111000010101010101101001011110111000100110101001010110000100000011101111111000000001000000000011000101010000000100100001010001100110100000001101011111110011110000001101101111110110000001001001100000111101100000011},
{784'b0111101100111110010010011100111001101100000111111000111000100110110011111110101111111010011000001010010111110011111001100000000111000000011100110110000010110101111011111010000000000010111111110011101100000000100000111111111001001100011011001111100010111010111100000101110110011001111011001001111101100000011000011110000010000001001111000010110101000110000101010100111000101101010100001000101101001000100111100010000000011100101101110100100000000011011000111111111101000001010101000000111111011000000011100101000000101111011010001100010000101000010101011111111101101111011110011111111110111010111101000111011101111100011111110011000011101111100010010000101000111111101110101010000001000110001110110111101000000001000011001010000110111111011000011011100111010100000100101101100001001100},
{784'b0010100000000011001100100010111001010000100001110011100111110111111000101111000101001000001101010100011011001101100010101100000001011000111111100000011100001101110000001000010111110100111110100001011111111110000111000111000010111111111100011111010111101010011111100001111111000001111100000100000111110011100011100100100000111100001001011100000000000111111111010010001010000000111111111110111110100000001111111111111000110110000011111111111101100101000010111111111111110101111111010111111111111100000110111110011111111110100100000111000100011111110000000001101011100010001101000000100010111100110100000000000000010101110111100000001000000101010110100110000000001000001110110011111000010000000010010001001010000000001001001001001111010100001011101000011011000101000011001011001010011110},
{784'b1010111001101101011010001000101000100001100000000111110001010000110000101001001001010111000111000110001000110111001111001001010111111111000010111110110011110110110001000000011110011110001111101001000010011101111010001000010100100110001111010000101101101001010001010000110010011110011011010110000010010011101000110000100000001101010110000011000010111000010100100100111001010111100000000010000001000111111110000101111000010101110111111001011111011110000001111101100101111111111001010111100100011111111111110001101110000100110111111100100111100001101001001111011000011111000100000110001111010000001000001001000010111001101110001000100010000010110001010100011000000000001110110000001000100011110001111011001000001101100101011001000111000110000101000001001000001010100011101000111101000000},
{784'b0011111001010011000101011111011110001100010011100010000100010101101110011001111100100011111111110001111111111010101011001111011101101110010001110010000001110010000001010100001000011100111111000110000100111000000111010111010101111110110000011111111001100110101111000011101000010001000110001000010110000001101001101001100001111100111111010101011100100111110010111001000001101010111111111101100001101111110001111111111110001011001110111100010011000000000010111111110011011010100101101111101000101110001000000110001110110011011011000001000100000001100001000001000010110100110000101000100011000110000100110011001000001001010101000010001101000010000101000010101010110000000000110111011101000000010101011110111011111111111000010111011110000001111111111110111101011101000000110111111100000000},
{784'b1000000000100011010100111101011100111000111010001000010110011011101010111001111100010011110001010000000000010000100111100000100000001101000101110000111110111000010110011110000111111111001000110110100000000111111011100010101100100011110011111100001110011001011011010111110000011101110010100010111110000111111110010110010111100000010001000001111000000100000000101001111101001010000000001101000001000000101000000001001101000000100000100000011001011000001000000010000001000110101111000100010000000110110001111110000101011010001110000100010010000111110001001101011110100000111111011111100010001000010111111000110000010110101010111111011111110011100110100111111111111101010100010110110010100011001110101111101011001000011010101111100101010001111110110100001010011000101110001111101001100111},
{784'b1011000110111110111000101101101000001011001110111101011101011100110000100000000100111011001001100000001101001101011101000000000011011111111010000110000001001011111100000100000101000000011111111001100010101000000001111111110000011010000000001111111110101111010100000011101111110001101110000001110111100100110001101001001110110000000000011110000011111001001010000101110100001000111100011110011011010000000001100001101001101010111011011100011110001100001101001111000111100000011010000010110000111110000001110110010010001111110000011111000111110100011110000000000011101101000111111000001110011011110011111100000001010010111100111110111000010111100101011101111010000000010001011101110000000000010111000110111011011000000000000011110001100111001000000000110001010011110111110111111010011011},
{784'b0111100011100110100101000101000000100000001000011001110010010010100110101011101010110000001111111111110110010010001101011111111111110110110100100011011111111111101010101100011010111111111011100111011011111110101111100100110001111010111001100000000001011111101111001000000010000011010011111000000000100000000011000010000010111111000000000111110000110111111100000001000000000001011111110000001101001000000000111110100000010110000000000111110010010001000000000000010100110010110001111000000000010101110110100001110000000010001111111010001111100000000111111111110110101111111011101110111100111010111111111111111111111100011111111111111101111111101001001111111111111101111110011000001111111101001010100101000001110111111000101010010100110101111011101111100101010011000011001011010101010100},
{784'b1010100110010001100010010010001101010100011110110010100001100010110011101011001011011010110000010100001110101110010100100001110001000100011101110011010000101100101001010000100101000000000100110011100101011111000101110001011000111011110011001111001110000000111111111100100111110101010011110111111010111111000000101111111111100011111110111011011111111110110111111011000011111111100101111111000110111111110000001101011100100100001111011010001011010100000001011111000101100000010111000000010101000011010000110110000000000000110000001011101101100000001111011010001101000001001011111110100000001100000001011111000111110010100000001111111110000001110000100011111111111100010000011110100011111111111010000111011111000111111010001100001000000001001100101101000011000110001001101000011101011001},
{784'b1111101111111100110010101100111011011001011011011001111110010111010011111111000101011101011101111111001101011110111011001110001111000111011010101010010011101000101001000110000011001010010011010111111000001000000000000101110110110101111110000011001110111111010100111000001111100011110111010111100011111100011110000111111111111011000110101110011001011111100000011010001011100000011110000000001110000000000101110101010011011011000000010010000000000110101100000111100010110001001001010100001111001111110100110111100000111000101111010110000000000001100011100011001111000000001111001011101101001101000000001110110010111110111000000000111010101111111011010000000001010000111011011001101001000011101010111010100111001001100110001100101010110111011001100001111001101110110101111110010110111111},
{784'b0000001010110011000000010000000011010000100000001110000010000101001111010001000000110000000100111110101000001000100010100111111110111100000110111010111111011011011011001111001111111100011111000100001001011111100111101000001100101111111100000110000000010001100111110000110000000100001001111110000001011000000001000111111000001111111000000001000111000000111111111110000001111100000001111111111000000001110100001111111101100101010111111100011111111001100000111111100011111111110101000101000000001111110111101011101111101111111111111100000100101101001101111111011010011111001011010011110110010010011010001100101111100100101101000111111110111110101000000010010011110010011000110001101101011011010001000000100010111011111100110001110010110000000110110000101000000010001100001001100000010001},
{784'b0010011111110011011011011111111111101101111001000101111010010111000100101101010110011011101100000000001000101010010110000000000000000010111000000010010000000000000000001100011000010010000000011010100111111010111110101101011101110100111010111111110111011010010100011111111110101111110111010111011110111011111100111111111000000110000011111001111111100000000000001111111011111111100000000100011101100111111101001111101010010111001111111011110111010001111110011111111011001011001001101000111111111101010010001111100000000101000100101001011100000000000011000000000011100000000000000111000111011110000000000110101011110101010100000001101000000011000100011001111000000100010101101111110100111011101011111011110100100001001101100111110111011111100100111010001100111000110001111001011101010100},
{784'b0101111100111001010101010101110000111100101001001000110001110100110100111011011101110001001000100000010101010101111111100001000000111011100111010010110000000111111110110000001111010000011111110111000000001110100001111110101010010001101111000011111001111011101111111000011111100011011001111111100001111110000010101110111000001111110000110111010000000001111111101110001111010000011011111100001010111100101011111111100010111101100100110111111100000101110111011000001111110000001101011000000111110100000001101111100000010001100000000110101111010000000010000000101001011010000000001100000000001101010111100000100100111100110001101000110011111100101100111001000000011111110111011111011111100000010011111101100001111110100000110110011110110101011100111011001110011111010101110001000000111011},
{784'b1010111110011111110101011011010010111100011010101011010011000001111110011001111000001011100110111110111111110101011001100011010101111111100000101010110000010100100110011011101000000000010000000001110010000101100001000000011101001101000100000000000000011110000000101111000000000000010011011101110001110000000110100000001111001111100000001101000111111101111110100111011111110011100011111100111111000101111110011111100010011100101111110001111110011011111111111111001111111110011110011111111110111111011111001111000011111011111101101110111111000001111111110101110100101000000000001001000001100001000000000000000000011000011100000000000000000000001010010000000000000000001000111110110001100000000011011110110011101101101111001011000011001101001000011110100111111111001111111110110110101111},
{784'b1110111011001001111100011111011010011000010011110101100101111010110000111111110111010111011010110110111110110000001101111000010101100001111001111110000001011110000000100011111110000011111000000111001010011000011111000000001010101111100001111100000010001110111110000111100000101001101111010000111100000010110011100000000111110000011000010110010101111110001011110001101101101111111111001010001111110000111111101010001100010101100001111101110011101000100100000001000011110110010101100000000000001110001100000111000000000001100011010001100010000000111000100100001010011010000001100110010011011111101111101110101110001110010111111111111000110100110110101101011111100001100011101001101111111010011001110011001010101101111101000110111111111001001011010011111011110010111111111001001011101110},
{784'b0001001110001000110101101110011110011100010110111010101110111101011100000011011010101100101110001100110000110000101011111010110000001010011010101101000000110100110000111010110000001110000011000001010111000001000000010111000000111110011001010001110100110110000000100101101111100000000110011000000010010010001100000010000000010000101000101110100001011110000101111111001001001010111111110011111011110111001010111010110011010001111000001100100111101110001001011100101101111001010001000111010111111110100011111111101000001111001010110011101100010000111111111110010110001101011110011110111010111111110011100001111100111101101000110111001100011111100110111110010001011101000100000110110001010001000011100101101000100000000000010111101101001100010100001010011010101111101010111100001011101110},
{784'b1010000100001001001000110100100000001010100110110000001101110001111111001111010110000001101111111101100100111100101011100101011000000001010100011010011101110000011111101100000000000111001011011111001010000001111111001100011000010100000001111100101110000110000000111110011000010001000001010111111001110001000111110011011000101010101100110010011010000010010011011100000100000100000000000110110000100111000001001000100111001101001100000010000000000100011010111111001100000000000001110111111111110000001001101110100111111111110100010111000000111111111110110001001100000001101110100110010010101100001111111110111011110110000111100111110000000001000011100001011000000111101110111010000000000000010111001111100110000000000101001110111100001101101111111110011101101000111111110010010001011011},
{784'b1111011101101100110010010001110101100111110111110110111111101001111000001010110111101111111100001001000000110010100100101101000000111110110110111110101010111100111101101100111010011111111001010001101001001110010111110100101110101000000100100011110000111110000000111101111110000000110101010011100111111000001110010011111101011111100000011110011111101011111111100111000011111101110111111000011001001011100011111110000011101110000000000111110000000110100001010001111111000001001111111000100110110100000001001011100001110110000001100111111110001001000000001010010001000000100000000100110110001110010010001000100101001100111100010010001000000011011001011101000001100000000100110010001000010011000111110001111111000100001011111000110110011111110101010011101011011101111100101110000011111111},
{784'b1101001100000111101100101010100001100001001000101011100100011010010110011111100100010111100010111101101100000100001000111111111010001010001101101111111111010000000000010101001111111100000010000100000111111111100000000000010100011111111100000001001001010011111111100000010101100111011011111110000111111100111101001010110000011111101101000000100111100011111101100010010011000011000100111100010010011110000000011111101101100111001110000001010111111010000000110000000111111011100110101001000001111111000110010000100000000111111110100011010110100000111111100001011000101011000011111110100010010011000010001111111100011000011100000000010011001001101010001011000001011110011000101011011101000000111100011000111111011111000011001010000100100000001010000001100100001010000000010110110101111011}};

logic signed  [63:0][127:0] l1_weights = 
{{128'b11001011101110011001110110110101100010110011110101101101010010001110011111000011111100111000011100000111011010111001000010101011},
{128'b01110111100101110110100110101011101011001010010110011111001110100010111001101100001010011101000101011011101010010100110111000011},
{128'b11001011000011111001100110000010001110100101101110111111100010110111000000000100110000001000010101110111000111010011011101000010},
{128'b10111100111010011000110001010111010011011001111101110000011010011011001110000010100100100111000010100101011000111101001100111001},
{128'b11011110001010111000000110100101001001111011101010101111100000010010111000010001101100001001010101100101011100100011001101111010},
{128'b01100010000111001001000111101001001101100011000110100111011100101010100011000101110011011110110001001000110011110101011001110100},
{128'b11001101100011000001100010101101011101000001101110000111010111001011101011010101110111101110101000001110100101110001011101001110},
{128'b01000001010101000011011011000100111110111110100101110011101100010100000100111110100111110001101010000100000111100111001100001101},
{128'b00101010101101101101110001100011011011101100010111011011001010011010101100000111101010011001011101011101111010010100101000011001},
{128'b00010110101100001001111001110001100010111010010101111100001001010010011111011010110101110011001101101101010110011001100011100001},
{128'b01111110110110011010010010101000000011110101111001001100110000101000111101001101100110011100010010010101111011110100111101011110},
{128'b01100110000011111110100000101101010001001000111111010010000101100010111001101100000110110001100001011000110000000100011000000001},
{128'b11011010000100111110100100110001000010101000011110101001111101110000011011001011101100010110100111110101000110010010011110011001},
{128'b00010101011111000111001101001100010100011110100010100000110101011010001000110111100001110111001011001000100000101011010001011100},
{128'b10011010100000101110110110100011100011101110011101110101110001100100110011001001000110011001100010110000000111011101101110000000},
{128'b01111101011101110110101111001100010011111100100100011001001000111100000111110010011001000011100111101011100000001000110111111001},
{128'b00101010000010001010001011101000011001111101011001010110011010101000100110001101110011011000010111001101111011011110111010000100},
{128'b01110111110100111110110010101110100010111010001010010101101111100110101000101001001111011100110001000101001011000100010101110111},
{128'b11110110111111101000100011100101000000111111010011101001100000011111101101000001001010011110110011111001011010000110000011010001},
{128'b00000011101110110110110001111000100010111000010001000100000011000010101111111011100000010011000000111111011010111000100010111001},
{128'b10001110100011110001000011110000010111100001000100100011010111011011100010010000110011101010101010101100110100011001111100101001},
{128'b00000101100001000110110110001101100101000010001110001010110011100011001001101100001001101100100100011010100101101101001101000101},
{128'b01101110100100001000110110100110000010101111011011011100001100101010101001101101100110010101011100001111110011110100001010000101},
{128'b01011011001000110001011010110010101101110000101101111111101000101110000011011100110001001100011000100011001111111100101100101110},
{128'b01101000000101001001000111101001001100111011000111100011111110101011000011011101110011011110110111001000110110010100011000100010},
{128'b00010101011001010011010110101000011001110010000101100001101100011011000110110000100001010111010011100000010000011101110001111000},
{128'b01110011111101100111100100001110110011111010000010101001000110010010011001010000101000000111010101000101100010100101000011011011},
{128'b00110010000010010000011011011000001001111110001001101000111110101101010110001111100011011010010010010001011111001110110000111100},
{128'b11101000010010011000001001010000011100111101010011101010110110111101110100111110000011111010011011111000110101001010011010110100},
{128'b11100100000101111101011111110011101110101110000111101011101110111001010011111101010011011111000111010010110110110101010010000010},
{128'b01111101010110011000010111111011100001000010101010000011000001111001111001101101111100001101000111010101110000100111000000111100},
{128'b01100100100101000001011011001110111000000100010011001010000110000001110101000111010101111000011001011000110000100111111010000100},
{128'b10000111100110101110111011010010100000110110111001011101001011000000100011111111011111011001101000011111111011110110101010000101},
{128'b11101000110111010010110110100101011011100101100110111011110100111011111110010001111010101100111111101001110110100000011000010011},
{128'b00101010001110111011011111000011011101100001100111011011010110011000010011000111111010011100110011010101110110110010001000011100},
{128'b10111100010000010010100100000110010110011111001010101100011111111100101100100110001101000000000111100110100001001100010101110101},
{128'b01101101000101101101011110101001100111100011000100111111101010101101100011011101011001011100111111000010010111011101011011100010},
{128'b10001000000101111100101101000001111001001100010101111110010000010100000100011110100010010001001100011111011100110010111110000001},
{128'b01101100101000111011011010001010010101110110100101111110111000011100010111001101110101011100010001000110111011111110011000001010},
{128'b01111110110100110110111100010110101001111110000000011101101000101100111100100000101100000001011110010111001011001110000101111101},
{128'b11110110011101011101011111111001100000111011000011101001101110111101010101101011001011011111111001010000110110000111000011110011},
{128'b10001001000001000111100110001101100111000101101110111011110110110101111010000100011001100110101110100110010101110011011101101110},
{128'b00110010011101001100111101110101110000011010110010000000000000011011111100110010100010110111001101011001110000101101100011011001},
{128'b00011101100011000011100000000110000101000000111110110100010001000010101010000101111111100101101000001111101000110000101101001000},
{128'b11011010110010011000100100000111011001100001011110111110110110011110011001100111101010101000010110100101101100111111011101011110},
{128'b00101100000101000000110001000100010011001110000101010000101000101100000000011010000011010001100111010010111000011100010111000001},
{128'b01010011111110011011110010100110000010111010100000000100111110001010001110010001110100110101100000110100001010110101110101111111},
{128'b10000111011010000000000001111101110001010001011001100000010101000011001011011101010110101010001010111001100101100111101000000100},
{128'b00110100000010100010001000011000010101010100001000011001101011100101100010111110011101000100011001010010011111001110100000011110},
{128'b11001001001101011111100110110101000011100110001100111101101110100011000011011101000101100111101101110011000111010011101010001010},
{128'b01011101011101010101100100110101111110000011100110001001000011111101001100010000001101101110101111110100000101000111010101111011},
{128'b00110100000110110110001010000100010000111010000001000100101010100100001101110011010001010001101100111011000011011110100111111101},
{128'b01110101111001010111001101001110011101110111000011010110011101111110101110110100111011100000100011000010111000001100010101110000},
{128'b10010011101000110110011001010010100101110110011001011000001001000101010101101111000001001000010110110011001111001110100110100100},
{128'b11101010010111011001001111000000011110101101001010111011110010000110110010111101101011011010010111101101110110011000011000000010},
{128'b00111100111000111010110010000010001111111111000100011001101110111100110110100001101100000111010011010111001010001100011101111111},
{128'b10000001011101101101101001010001100111001111001000010011000011110111110110100010001000100111101111111101010100001011000010101011},
{128'b01110110011111101000001011111001010000011011011011100001101100101011111001100011010010011111110011011000100110001111000010111000},
{128'b00100100001101110110100101110000111000001000010101111000110011001010100100100000000110010001001001001000110001110100101110000011},
{128'b11111100011101011011000001011111010001011110101011101011110001110111110010100110000111100110101111111000110101001011010010110000},
{128'b00101000000101010101000111101110010101000111100110010010111100111101100000100101000111010111111101010000110000010101011000001101},
{128'b11001000110101110110100100110111111111100000111010011110101011101101110101101100000010101000011110111001100111101011011110000001},
{128'b01101010000111101101111111110001011010101010010101111001111010001010000110111001110010010010100001001101111010111000110011011011},
{128'b10000111110010101011000000101100101100110011001000000101100001001110101011010101110100011100011000100000001001110001001001111110}};

logic [9:0][63:0] out_weights =
{{8'b1011110010101000100000010011101001111111010010001010111100000100},
{8'b1110111010110100011001000010001101100001101110110010000001000101},
{8'b1011101001001010000111010000000000000100010110110110010010000101},
{8'b1111100010111011111100100010000001010101001111100011000100100110},
{8'b1011111011001110001010001010011001101000111010100110001111011010},
{8'b1001000011110010101110100001111111100100101000010000011011100110},
{8'b0011111010111010111010101101101001110010000110110000101001010001},
{8'b0111100000011010011001000010111001011001110110001110011111010100},
{8'b1110111010111010100011111000010111101110010111000100001000101110},
{8'b1010110011101010111100111111011010101011100010100101011101000011}};